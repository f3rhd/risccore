module control_unit(
    input logic[31:0] instr,
    output logic[25:0] ctrl_signals
);
    // # INPUT = OP(7)+FUNC(3)+FUNC(7)mm_type_select(3) + r
    //output = j(1) + beq(1) + bne(1) + blt(1) + bge(1) + bltu(1) + bgeu(1) + + imm_type(3) + REG_WRITE(1) + ALU_B_OPERAND_SELECT(1) + ALU_CMP_TYPE(1) + ALU_OP_TYPE(4) + RAM_READ_TYPE(3) + RAM_WRITE_TYPE(2) + WRITE_DATA_SELECT(3) + PC_SELECT_B_OPERAND_SELECT(1)
    always_comb begin
        logic[16:0] pla_input;
        pla_input[16:10] = instr[6:0];
        pla_input[9:7] = instr[14:12];
        pla_input[6:0] = instr[31:25];

        casez(pla_input)
            17'b0000011_000_??????? : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_1_0_0010_101_00_101_0;
            17'b0000011_001_??????? : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_1_0_0010_011_00_101_0;
            17'b0000011_010_??????? : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_1_0_0010_001_00_101_0;
            17'b0000011_100_??????? : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_1_0_0010_100_00_101_0;
            17'b0000011_101_??????? : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_1_0_0010_010_00_101_0;
            17'b0010011_000_??????? : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_1_0_0010_000_00_011_0;
            17'b0010011_001_0000000 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_1_0_0011_000_00_011_0;
            17'b0010011_010_??????? : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_1_0_0011_000_00_010_0;
            17'b0010011_011_??????? : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_1_1_0011_000_00_010_0;
            17'b0010011_100_??????? : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_1_0_0101_000_00_011_0;
            17'b0010011_101_0000000 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_1_0_0100_000_00_011_0;
            17'b0010011_101_0100000 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_1_0_0101_000_00_011_0;
            17'b0010011_110_??????? : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_1_0_0111_000_00_011_0;
            17'b0010011_111_??????? : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_1_0_0001_000_00_011_0;
            17'b0010111_???_??????? : ctrl_signals =  26'b0_0_0_0_0_0_0_010_1_0_0_0000_000_00_111_0;
            17'b0100011_000_??????? : ctrl_signals =  26'b0_0_0_0_0_0_0_100_0_1_0_0010_000_10_000_0;
            17'b0100011_001_??????? : ctrl_signals =  26'b0_0_0_0_0_0_0_100_0_1_0_0010_000_01_000_0;
            17'b0100011_010_??????? : ctrl_signals =  26'b0_0_0_0_0_0_0_100_0_1_0_0010_000_11_000_0;
            17'b0110011_000_0000000 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_0010_000_00_011_0;
            17'b0110011_000_0100000 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_0110_000_00_011_0;
            17'b0110011_001_0000000 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_0011_000_00_011_0;
            17'b0110011_010_0000000 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_0000_000_00_010_0;
            17'b0110011_011_0000000 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_1_0000_000_00_010_0;
            17'b0110011_100_0000000 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_0000_000_00_011_0;
            17'b0110011_101_0000000 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_0100_000_00_011_0;
            17'b0110011_101_0100000 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_0101_000_00_011_0;
            17'b0110011_110_0000000 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_0111_000_00_011_0;
            17'b0110011_111_0000000 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_0001_000_00_011_0;
            17'b0110111_???_??????? : ctrl_signals =  26'b0_0_0_0_0_0_0_010_1_0_0_0000_000_00_100_0;
            17'b1100011_000_??????? : ctrl_signals =  26'b0_1_0_0_0_0_0_111_0_0_0_0000_000_00_000_0;
            17'b1100011_001_??????? : ctrl_signals =  26'b0_0_1_0_0_0_0_111_0_0_0_0000_000_00_000_0;
            17'b1100011_100_??????? : ctrl_signals =  26'b0_0_0_1_0_0_0_111_0_0_0_0000_000_00_000_0;
            17'b1100011_101_??????? : ctrl_signals =  26'b0_0_0_0_1_0_0_111_0_0_0_0000_000_00_000_0;
            17'b1100011_110_??????? : ctrl_signals =  26'b0_0_0_0_0_1_0_111_0_0_1_0000_000_00_000_0;
            17'b1100011_111_??????? : ctrl_signals =  26'b0_0_0_0_0_0_1_111_0_0_1_0000_000_00_000_0;
            17'b1100111_000_??????? : ctrl_signals =  26'b1_0_0_0_0_0_0_000_1_1_0_0010_000_00_110_1;
            17'b1101111_???_??????? : ctrl_signals =  26'b1_0_0_0_0_0_0_001_1_1_0_0000_000_00_110_0;
            17'b0110011_000_0000001 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_1000_000_00_011_0;
            17'b0110011_100_0000001 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_1001_000_00_011_0;
            17'b0110011_101_0000001 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_1010_000_00_011_0;
            17'b0110011_110_0000001 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_1011_000_00_011_0;
            17'b0110011_111_0000001 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_1100_000_00_011_0;
            17'b0110011_001_0000001 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_1101_000_00_011_0;
            17'b0110011_010_0000001 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_1110_000_00_011_0;
            17'b0110011_011_0000001 : ctrl_signals =  26'b0_0_0_0_0_0_0_000_1_0_0_1111_000_00_011_0;
            default:
                ctrl_signals = 26'd0;
        endcase
    end
endmodule








