module control_unit(
    input logic[31:0] instr,
    output logic[25:0] ctrl_signals
);
    // # INPUT = OP(7)+FUNC(3)+FUNC(7)mm_type_select(3) + r
    //output = j(1) + beq(1) + bne(1) + blt(1) + bge(1) + bltu(1) + bgeu(1) iEG_WRITE(1) + ALU_B_OPERAND_SELECT(1) + ALU_CMP_TYPE(1) + ALU_OP_TYPE(4) + RAM_READ_TYPE(3) + RAM_WRITE_TYPE(2) + WRITE_DATA_SELECT(3)
    always_comb begin
        logic[16:0] pla_input;
        pla_input[16:10] = instr[6:0];
        pla_input[9:7] = instr[14:12];
        pla_input[6:0] = instr[31:25];

        casez(pla_input)
            17'b0000011000??????? : ctrl_signals =  26'b00000000001100010101001010;
            17'b0000011001??????? : ctrl_signals =  26'b00000000001100010011001010;
            17'b0000011010??????? : ctrl_signals =  26'b00000000001100010001001010;
            17'b0000011100??????? : ctrl_signals =  26'b00000000001100010100001010;
            17'b0000011101??????? : ctrl_signals =  26'b00000000001100010010001010;
            17'b0010011000??????? : ctrl_signals =  26'b00000000001100010000000110;
            17'b00100110010000000 : ctrl_signals =  26'b00000000001100011000000110;
            17'b0010011010??????? : ctrl_signals =  26'b00000000001100011000000100;
            17'b0010011011??????? : ctrl_signals =  26'b00000000001110011000000100;
            17'b0010011100??????? : ctrl_signals =  26'b00000000001100101000000110;
            17'b00100111010000000 : ctrl_signals =  26'b00000000001100100000000110;
            17'b00100111010100000 : ctrl_signals =  26'b00000000001100101000000110;
            17'b0010011110??????? : ctrl_signals =  26'b00000000001100111000000110;
            17'b0010011111??????? : ctrl_signals =  26'b00000000001100001000000110;
            17'b0010111?????????? : ctrl_signals =  26'b00000000101000000000001110;
            17'b0100011000??????? : ctrl_signals =  26'b00000001000100010000100000;
            17'b0100011001??????? : ctrl_signals =  26'b00000001000100010000010000;
            17'b0100011010??????? : ctrl_signals =  26'b00000001000100010000110000;
            17'b01100110000000000 : ctrl_signals =  26'b00000000001000010000000110;
            17'b01100110000100000 : ctrl_signals =  26'b00000000001000110000000110;
            17'b01100110010000000 : ctrl_signals =  26'b00000000001000011000000110;
            17'b01100110100000000 : ctrl_signals =  26'b00000000001000000000000100;
            17'b01100110110000000 : ctrl_signals =  26'b00000000001010000000000100;
            17'b01100111000000000 : ctrl_signals =  26'b00000000001000000000000110;
            17'b01100111010000000 : ctrl_signals =  26'b00000000001000100000000110;
            17'b01100111010100000 : ctrl_signals =  26'b00000000001000101000000110;
            17'b01100111100000000 : ctrl_signals =  26'b00000000001000111000000110;
            17'b01100111110000000 : ctrl_signals =  26'b00000000001000001000000110;
            17'b0110111?????????? : ctrl_signals =  26'b00000000101000000000001000;
            17'b1100011000??????? : ctrl_signals =  26'b01000001110000000000000000;
            17'b1100011001??????? : ctrl_signals =  26'b00100001110000000000000000;
            17'b1100011100??????? : ctrl_signals =  26'b00010001110000000000000000;
            17'b1100011101??????? : ctrl_signals =  26'b00001001110000000000000000;
            17'b1100011110??????? : ctrl_signals =  26'b00000101110010000000000000;
            17'b1100011111??????? : ctrl_signals =  26'b00000011110010000000000000;
            17'b1100111000??????? : ctrl_signals =  26'b1_0_0_0_0_0_0_000_1100010000001101;
            17'b1101111?????????? : ctrl_signals =  26'b1_0_0_0_0_0_0_001_1100000000001100;
            17'b01100110000000001 : ctrl_signals =  26'b00000000001001000000000110;
            17'b01100111000000001 : ctrl_signals =  26'b00000000001001001000000110;
            17'b01100111010000001 : ctrl_signals =  26'b00000000001001010000000110;
            17'b01100111100000001 : ctrl_signals =  26'b00000000001001011000000110;
            17'b01100111110000001 : ctrl_signals =  26'b00000000001001100000000110;
            default:
                ctrl_signals = 26'd0;
        endcase
    end
endmodule








