module control_unit(
    input logic[31:0] instr,
    output logic[24:0] ctrl_signals
);
    // # INPUT = OP(7)+FUNC(3)+FUNC(7)mm_type_select(3) + r
    //output = j(1) + beq(1) + bne(1) + blt(1) + bge(1) + bltu(1) + bgeu(1) iEG_WRITE(1) + ALU_B_OPERAND_SELECT(1) + ALU_CMP_TYPE(1) + ALU_OP_TYPE(4) + RAM_READ_TYPE(3) + RAM_WRITE_TYPE(2) + WRITE_DATA_SELECT(3)
    always_comb begin
        logic[16:0] pla_input;
        pla_input[16:10] = instr[6:0];
        pla_input[9:7] = instr[14:12];
        pla_input[6:0] = instr[31:25];

        casez(pla_input)
            17'b0000011000??????? : ctrl_signals =  25'b0000000000110001010100101;
            17'b0000011001??????? : ctrl_signals =  25'b0000000000110001001100101;
            17'b0000011010??????? : ctrl_signals =  25'b0000000000110001000100101;
            17'b0000011100??????? : ctrl_signals =  25'b0000000000110001010000101;
            17'b0000011101??????? : ctrl_signals =  25'b0000000000110001001000101;
            17'b0010011000??????? : ctrl_signals =  25'b0000000000110001000000011;
            17'b00100110010000000 : ctrl_signals =  25'b0000000000110001100000011;
            17'b0010011010??????? : ctrl_signals =  25'b0000000000110001100000010;
            17'b0010011011??????? : ctrl_signals =  25'b0000000000111001100000010;
            17'b0010011100??????? : ctrl_signals =  25'b0000000000110010100000011;
            17'b00100111010000000 : ctrl_signals =  25'b0000000000110010000000011;
            17'b00100111010100000 : ctrl_signals =  25'b0000000000110010100000011;
            17'b0010011110??????? : ctrl_signals =  25'b0000000000110011100000011;
            17'b0010011111??????? : ctrl_signals =  25'b0000000000110000100000011;
            17'b0010111?????????? : ctrl_signals =  25'b0000000010100000000000111;
            17'b0100011000??????? : ctrl_signals =  25'b0000000100010001000010000;
            17'b0100011001??????? : ctrl_signals =  25'b0000000100010001000001000;
            17'b0100011010??????? : ctrl_signals =  25'b0000000100010001000011000;
            17'b01100110000000000 : ctrl_signals =  25'b0000000000100001000000011;
            17'b01100110000100000 : ctrl_signals =  25'b0000000000100011000000011;
            17'b01100110010000000 : ctrl_signals =  25'b0000000000100001100000011;
            17'b01100110100000000 : ctrl_signals =  25'b0000000000100000000000010;
            17'b01100110110000000 : ctrl_signals =  25'b0000000000101000000000010;
            17'b01100111000000000 : ctrl_signals =  25'b0000000000100000000000011;
            17'b01100111010000000 : ctrl_signals =  25'b0000000000100010000000011;
            17'b01100111010100000 : ctrl_signals =  25'b0000000000100010100000011;
            17'b01100111100000000 : ctrl_signals =  25'b0000000000100011100000011;
            17'b01100111110000000 : ctrl_signals =  25'b0000000000100000100000011;
            17'b0110111?????????? : ctrl_signals =  25'b0000000010100000000000100;
            17'b1100011000??????? : ctrl_signals =  25'b0100000111000000000000000;
            17'b1100011001??????? : ctrl_signals =  25'b0010000111000000000000000;
            17'b1100011100??????? : ctrl_signals =  25'b0001000111000000000000000;
            17'b1100011101??????? : ctrl_signals =  25'b0000100111000000000000000;
            17'b1100011110??????? : ctrl_signals =  25'b0000010111001000000000000;
            17'b1100011111??????? : ctrl_signals =  25'b0000001111001000000000000;
            17'b1100111?????????? : ctrl_signals =  25'b1000000000110001000000110;
            17'b1101111?????????? : ctrl_signals =  25'b1000000001110000000000110;
            17'b01100110000000001 : ctrl_signals =  25'b0000000000100100000000011;
            17'b01100111000000001 : ctrl_signals =  25'b0000000000100100100000011;
            17'b01100111010000001 : ctrl_signals =  25'b0000000000100101000000011;
            17'b01100111100000001 : ctrl_signals =  25'b0000000000100101100000011;
            17'b01100111110000001 : ctrl_signals =  25'b0000000000100110000000011;
            default:
                ctrl_signals = 25'd0;
        endcase
    end
endmodule








